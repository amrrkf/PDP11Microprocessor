library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

Entity rom is
port (
clk : in std_logic;
uAR : in std_logic_vector(7 downto 0);
CW : out std_logic_vector(31 downto 0) );
end entity rom;

architecture rom_arch of rom is
	type rom_type is array(0 to 255) of std_logic_vector(31 downto 0);

	signal rom : rom_type := (
0   =>  "00000001000101101000001011100000",
1   =>  "00000010001100100000000000000000",
2   =>  "00000011001001000000000000000000",
3   =>  "00000000000000000000000000000001",
4	=>	"00000000000000000000000110000000",
16	=>	"10111100100001100000001001011000",
17	=>	"10111100100001100000001000011000",
18	=>	"10111100100001100000010000111000",
20	=>	"00011101000000000000000000000000",
21	=>	"10111100100001100000101000011000",
22	=>	"10111100100001100000110000011000",
23	=>	"00011000000001100000000000000000",
24	=>	"00011001001100011000000000000000",
25	=>	"00011010100000000010000000000000",
26	=>	"00000000101000000000010000110000",
28	=>	"00000000100000000000100000010000",
29	=>	"00011110000001100000000000000000",
30	=>	"00011111001100011000000000000000",
31	=>	"00100000100000000010000000000000",
32	=>	"00100001000001100000111000000000",
33	=>	"00100010001100000010000000000000",
34	=>	"10111100101001100000100000011000",
35	=>	"00100100101100000010000000000000",
36	=>	"00100101000101100000001000000000",
37	=>	"00000000001100100000000000000000",
44	=>	"00010000000000000000000000001010",
46	=>	"11000000000000000000000000001110",
47	=>	"00110000000001100000000000000000",
48	=>	"00110001001100011000000000000000",
49	=>	"00110010011000000010000000000000",
50	=>	"00110011000001100000011000000000",
51	=>	"00110100001111001000000000000000",
52	=>	"00110101010000010000000100000000",
53	=>	"00110110000110000000000000000000",
54	=>	"00000000101000100000000000000000",
56	=>	"00111001010000100000000000000000",
57	=>	"00111010011000001010000010000000",
58	=>	"00111011000001100000000000100000",
59	=>	"00111100001010000000000000000000",
60	=>	"00000000001111000000000000000000",
65	=>	"10000001010000000100000000000010",
73	=>	"01001010010000001000000010000000",
74	=>	"01111010000000000000000000000000",
81	=>	"01010010010001101000001011100000",
82	=>	"01111000001110000000000000000100",
97	=>	"01100010010000000010000000000000",
98	=>	"01100011000001100000011000000000",
99	=>	"01100100001110001000000010000000",
100	=>	"01111000000000000000000000000100",
113	=>	"01110010000101101000001011100000",
114	=>	"01110011001100100000000000000000",
115	=>	"01110100001000000010000000000000",
116	=>	"01110101010001100000001000000000",
117	=>	"01110110001100001000000010000000",
118	=>	"01111000000000000000000000000100",
120	=>	"01111001001000001000000010000000",
121	=>	"01111010000000000000000000000000",
122	=>	"10000000001000000100000000000000",
128	=>	"10000001000000000000000000000010",
129	=>	"00101100010100000010000000001100",
137	=>	"10001010010100001000000010000000",
138	=>	"10111010000000000000000000000000",
145	=>	"10010010010101101000001011100000",
146	=>	"10111000001110100000000000000110",
161	=>	"10100010010100000010000000000000",
162	=>	"10100011000001100000011000000000",
163	=>	"10100100001110101000000010000000",
164	=>	"10111000000000000000000000000110",
177	=>	"10110010000101101000001011100000",
178	=>	"10110011001100100000000000000000",
179	=>	"10110100001000000010000000000000",
180	=>	"10110101010101100000001000000000",
181	=>	"10110110001100001000000010000000",
182	=>	"10111000000000000000000000000110",
184	=>	"10111001001000001000000010000000",
185	=>	"10111010000000000000000000000000",
186	=>	"00101100001000000010000000001100",
188	=>	"00000000001100010000000100000000",
189	=>	"00000000001110100000000000000000",
192	=>	"10111100000001100000000000111000",
195	=>	"10111100000001100000011000011000",
199	=>	"10111100000001100000111000011000",
200	=>	"10111100000001100001000000011000",
201	=>	"10111100000001100001001000011000",
202	=>	"10111100000001100001010000011000",
203	=>	"10111100000001100001011000011000",
204	=>	"10111100000001100001100000011000",
205	=>	"10111100000001100001101000011000",
206	=>	"10111100000001100001110000011000",
207	=>	"10111100000001100001111000011000",
211	=>	"10111100000001100000011000111000",
224	=>	"11100001000001100000000000000000",
225	=>	"00000000001100100000000000000000",
others => "00000000000000000000000000000000"
);
	begin
		process(clk) is
		  Begin
			if falling_edge(clk) then  
				CW <= rom(to_integer(unsigned(uAR)));
			end if;
		end process;

end architecture rom_arch;
